module hexdecoder
(
input [3:0] in,
output [6:0] out
);

assign out =
    (in == 5'h00) ? 7'b1000000 :
    (in == 5'h01) ? 7'b1111001 :
    (in == 5'h02) ? 7'b0100100 :
    (in == 5'h03) ? 7'b0110000 :
    (in == 5'h04) ? 7'b0011001 :
    (in == 5'h05) ? 7'b0010010 :
    (in == 5'h06) ? 7'b0000010 :
    (in == 5'h07) ? 7'b1111000 :
    (in == 5'h08) ? 7'b0000000 :
    (in == 5'h09) ? 7'b0010000 :
    (in == 5'h0A) ? 7'b0001000 :
    (in == 5'h0B) ? 7'b0000011 :
    (in == 5'h0C) ? 7'b1000110 :
    (in == 5'h0D) ? 7'b0100001 :
    (in == 5'h0E) ? 7'b0000110 : 
	 7'b0001110;
     
endmodule